module Instruction_Memory(
    input [31:0] address,
    output [31:0] data
);
    reg [31:0] mem [80:0];
    initial begin
// Initialize x1 = 0, x2 = 1
    mem[0] = 32'h00000093; // addi x1, x0, 0
    mem[1] = 32'h00100113; // addi x2, x0, 1

    // Store first two numbers to memory 0(x0) and 4(x0)
    mem[2] = 32'h00102023; // sw x1, 0(x0) = 0
    mem[3] = 32'h00202223; // sw x2, 4(x0) = 1

    // Generate Fibonacci numbers (fully unrolled, storing each result to memory)
    mem[4]  = 32'h002081B3; // add x3, x1, x2 => 0+1=1
    mem[5]  = 32'h00302423; // sw x3, 8(x0) => 1
    mem[6]  = 32'h002000B3; // add x1, x0, x2 => x1=1
    mem[7]  = 32'h00300133; // add x2, x0, x3 => x2=1

    mem[8]  = 32'h002081B3; // add x3, x1, x2 => 1+1=2
    mem[9]  = 32'h00302623; // sw x3, 12(x0) => 2
    mem[10] = 32'h002000B3; // add x1, x0, x2 => x1=1
    mem[11] = 32'h00300133; // add x2, x0, x3 => x2=2

    mem[12] = 32'h002081B3; // add x3, x1, x2 => 1+2=3
    mem[13] = 32'h00302823; // sw x3, 16(x0) => 3
    mem[14] = 32'h002000B3; // add x1, x0, x2 => x1=2
    mem[15] = 32'h00300133; // add x2, x0, x3 => x2=3

    mem[16] = 32'h002081B3; // add x3, x1, x2 => 2+3=5
    mem[17] = 32'h00302A23; // sw x3, 20(x0) => 5
    mem[18] = 32'h002000B3; // add x1, x0, x2 => x1=3
    mem[19] = 32'h00300133; // add x2, x0, x3 => x2=5

    mem[20] = 32'h002081B3; // add x3, x1, x2 => 3+5=8
    mem[21] = 32'h00302C23; // sw x3, 24(x0) => 8
    mem[22] = 32'h002000B3; // add x1, x0, x2 => x1=5
    mem[23] = 32'h00300133; // add x2, x0, x3 => x2=8

    mem[24] = 32'h002081B3; // add x3, x1, x2 => 5+8=13
    mem[25] = 32'h00302E23; // sw x3, 28(x0) => 13
    mem[26] = 32'h002000B3; // add x1, x0, x2 => x1=8
    mem[27] = 32'h00300133; // add x2, x0, x3 => x2=13

    mem[28] = 32'h002081B3; // add x3, x1, x2 => 8+13=21
    mem[29] = 32'h003020A3; // sw x3, 32(x0) => 21
    mem[30] = 32'h002000B3; // add x1, x0, x2 => x1=13
    mem[31] = 32'h00300133; // add x2, x0, x3 => x2=21

    mem[32] = 32'h002081B3; // add x3, x1, x2 => 13+21=34
    mem[33] = 32'h003022A3; // sw x3, 36(x0) => 34
    mem[34] = 32'h002000B3; // add x1, x0, x2 => x1=21
    mem[35] = 32'h00300133; // add x2, x0, x3 => x2=34

    mem[36] = 32'h002081B3; // add x3, x1, x2 => 21+34=55
    mem[37] = 32'h003024A3; // sw x3, 40(x0) => 55
    mem[38] = 32'h002000B3; // add x1, x0, x2 => x1=34
    mem[39] = 32'h00300133; // add x2, x0, x3 => x2=55

    mem[40] = 32'h002081B3; // add x3, x1, x2 => 34+55=89
    mem[41] = 32'h003026A3; // sw x3, 44(x0) => 89
    mem[42] = 32'h002000B3; // add x1, x0, x2 => x1=55
    mem[43] = 32'h00300133; // add x2, x0, x3 => x2=89

    mem[44] = 32'h002081B3; // add x3, x1, x2 => 55+89=144
    mem[45] = 32'h003028A3; // sw x3, 48(x0) => 144
    mem[46] = 32'h002000B3; // add x1, x0, x2 => x1=89
    mem[47] = 32'h00300133; // add x2, x0, x3 => x2=144

    mem[48] = 32'h002081B3; // add x3, x1, x2 => 89+144=233
    mem[49] = 32'h00302AA3; // sw x3, 52(x0) => 233
    mem[50] = 32'h002000B3; // add x1, x0, x2 => x1=144
    mem[51] = 32'h00300133; // add x2, x0, x3 => x2=233

    mem[52] = 32'h002081B3; // add x3, x1, x2 => 144+233=377
    mem[53] = 32'h00302CA3; // sw x3, 56(x0) => 377
    mem[54] = 32'h002000B3; // add x1, x0, x2 => x1=233
    mem[55] = 32'h00300133; // add x2, x0, x3 => x2=377

    mem[56] = 32'h002081B3; // add x3, x1, x2 => 233+377=610
    mem[57] = 32'h00302EA3; // sw x3, 60(x0) => 610
    mem[58] = 32'h002000B3; // add x1, x0, x2 => x1=377
    mem[59] = 32'h00300133; // add x2, x0, x3 => x2=610

    mem[60] = 32'h002081B3; // add x3, x1, x2 => 377+610=987
    mem[61] = 32'h00302023; // sw x3, 64(x0) => 987
    mem[62] = 32'h002000B3; // add x1, x0, x2 => x1=610
    mem[63] = 32'h00300133; // add x2, x0, x3 => x2=987

    mem[64] = 32'h002081B3; // add x3, x1, x2 => 610+987=1597
    mem[65] = 32'h00302223; // sw x3, 68(x0) => 1597
    mem[66] = 32'h002000B3; // add x1, x0, x2 => x1=987
    mem[67] = 32'h00300133; // add x2, x0, x3 => x2=1597

    mem[68] = 32'h002081B3; // add x3, x1, x2 => 987+1597=2584
    mem[69] = 32'h00302423; // sw x3, 72(x0) => 2584
    mem[70] = 32'h002000B3; // add x1, x0, x2 => x1=1597
    mem[71] = 32'h00300133; // add x2, x0, x3 => x2=2584

    mem[72] = 32'h002081B3; // add x3, x1, x2 => 1597+2584=4181
    mem[73] = 32'h00302623; // sw x3, 76(x0) => 4181
    mem[74] = 32'h002000B3; // add x1, x0, x2 => x1=2584
    mem[75] = 32'h00300133; // add x2, x0, x3 => x2=4181
    
    mem[76] = 32'h002081B3; // add x3, x1, x2 => 2584+4181=6765
    mem[77] = 32'h00302423; // sw x3, 80(x0) => 6765
    end
    
    assign data = mem[address[31:2]];
endmodule